
package fifo_pkg;
 `include"uvm_macros.svh"
	import uvm_pkg::*;

	int no_of_transactions = 200;

  //typedef uvm_config_db#(virtual io_if) vif_config;
  // typedef virtual fiof_if d_vif;
   //typedef virtual fiof_if im_vif;
  // typedef virtual fiof_if om_vif;
   
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/rtl/defines.v"	
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/input_agent/input_agent_config.sv"
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/input_agent/input_trans.sv"
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/input_agent/input_sequence.sv"
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/input_agent/input_sequencer.sv"
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/input_agent/input_driver.sv"
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/input_agent/input_monitor.sv"
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/input_agent/input_agent.sv"
  
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/output_agent/output_agent_config.sv"
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/output_agent/output_trans.sv"
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/output_agent/output_monitor.sv"
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/agents/output_agent/output_agent.sv"
   
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/tb/scoreboard.sv"
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/tb/env_config.sv"  
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/tb/env.sv"
  
  `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/test/test_top.sv"
   `include "/export/home/durga_b21/UVM/FIFO_uvm_durga/test/test_fifo.sv"
   

endpackage : fifo_pkg
